`timescale 1ns / 1ps


module encoder_8x3_dataflow_tb;
reg d0,d1,d2,d3,d4,d5,d6,d7;
wire a,b,c;
encoder_8x3_dataflow dut(.d0(d0),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.d5(d5),.d6(d6),.d7(d7),.a(a),.b(b),.c(c));
initial begin
/*d0=1; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0;
#10
d0=0; d1=1; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0;
#10
d0=0; d1=0; d2=1; d3=0; d4=0; d5=0; d6=0; d7=0;
#10
d0=0; d1=0; d2=0; d3=1; d4=0; d5=0; d6=0; d7=0;
#10
d0=0; d1=0; d2=0; d3=0; d4=1; d5=0; d6=0; d7=0;
#10
d0=0; d1=0; d2=0; d3=0; d4=0; d5=1; d6=0; d7=0;
#10
d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=1; d7=0;
#10
d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=1;*/
d0=8'b1000_0000;#10
d1=8'b0100_0000;#10
d2=8'b0010_0000;#10
d3=8'b0001_0000;#10
d4=8'b0000_1000;#10
d5=8'b0000_0100;#10
d6=8'b0000_0010;#10
d7=8'b0000_0001;#50

$finish;
end
endmodule
